module hello_world;

  initial begin
    $display("Hello, World!");
    $finish; // End simulation
  end

endmodule